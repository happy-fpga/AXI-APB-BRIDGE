VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO axi_apb_bridge
  CLASS BLOCK ;
  FOREIGN axi_apb_bridge ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1800.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.620 10.640 170.220 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 322.220 10.640 323.820 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.820 10.640 477.420 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 629.420 10.640 631.020 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 783.020 10.640 784.620 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.620 10.640 938.220 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1090.220 10.640 1091.820 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1243.820 10.640 1245.420 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1397.420 10.640 1399.020 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1551.020 10.640 1552.620 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.620 10.640 1706.220 1787.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.380 1794.700 21.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 173.560 1794.700 175.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.740 1794.700 328.340 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 479.920 1794.700 481.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 633.100 1794.700 634.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 786.280 1794.700 787.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 939.460 1794.700 941.060 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1092.640 1794.700 1094.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1245.820 1794.700 1247.420 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1399.000 1794.700 1400.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1552.180 1794.700 1553.780 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1705.360 1794.700 1706.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.320 10.640 166.920 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.920 10.640 320.520 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 472.520 10.640 474.120 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 626.120 10.640 627.720 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 779.720 10.640 781.320 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 933.320 10.640 934.920 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1086.920 10.640 1088.520 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1240.520 10.640 1242.120 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1394.120 10.640 1395.720 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1547.720 10.640 1549.320 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1701.320 10.640 1702.920 1787.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.080 1794.700 18.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 170.260 1794.700 171.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 323.440 1794.700 325.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 476.620 1794.700 478.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 629.800 1794.700 631.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 782.980 1794.700 784.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 936.160 1794.700 937.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1089.340 1794.700 1090.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1242.520 1794.700 1244.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1395.700 1794.700 1397.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1548.880 1794.700 1550.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1702.060 1794.700 1703.660 ;
    END
  END VPWR
  PIN apb_paddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END apb_paddr[0]
  PIN apb_paddr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 463.770 1796.000 464.050 1800.000 ;
    END
  END apb_paddr[10]
  PIN apb_paddr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END apb_paddr[11]
  PIN apb_paddr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1553.840 1800.000 1554.440 ;
    END
  END apb_paddr[12]
  PIN apb_paddr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1796.000 1346.330 1800.000 ;
    END
  END apb_paddr[13]
  PIN apb_paddr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END apb_paddr[14]
  PIN apb_paddr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END apb_paddr[15]
  PIN apb_paddr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 573.250 1796.000 573.530 1800.000 ;
    END
  END apb_paddr[16]
  PIN apb_paddr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1292.040 1800.000 1292.640 ;
    END
  END apb_paddr[17]
  PIN apb_paddr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 741.240 1800.000 741.840 ;
    END
  END apb_paddr[18]
  PIN apb_paddr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END apb_paddr[19]
  PIN apb_paddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END apb_paddr[1]
  PIN apb_paddr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 217.640 1800.000 218.240 ;
    END
  END apb_paddr[20]
  PIN apb_paddr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 363.840 1800.000 364.440 ;
    END
  END apb_paddr[21]
  PIN apb_paddr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1796.000 1401.070 1800.000 ;
    END
  END apb_paddr[22]
  PIN apb_paddr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END apb_paddr[23]
  PIN apb_paddr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END apb_paddr[24]
  PIN apb_paddr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END apb_paddr[25]
  PIN apb_paddr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 102.040 1800.000 102.640 ;
    END
  END apb_paddr[26]
  PIN apb_paddr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 537.240 1800.000 537.840 ;
    END
  END apb_paddr[27]
  PIN apb_paddr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END apb_paddr[28]
  PIN apb_paddr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1043.370 1796.000 1043.650 1800.000 ;
    END
  END apb_paddr[29]
  PIN apb_paddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1145.840 1800.000 1146.440 ;
    END
  END apb_paddr[2]
  PIN apb_paddr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1785.040 1800.000 1785.640 ;
    END
  END apb_paddr[30]
  PIN apb_paddr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END apb_paddr[31]
  PIN apb_paddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 1796.000 216.110 1800.000 ;
    END
  END apb_paddr[3]
  PIN apb_paddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1783.970 1796.000 1784.250 1800.000 ;
    END
  END apb_paddr[4]
  PIN apb_paddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1796.000 1153.130 1800.000 ;
    END
  END apb_paddr[5]
  PIN apb_paddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 602.230 1796.000 602.510 1800.000 ;
    END
  END apb_paddr[6]
  PIN apb_paddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END apb_paddr[7]
  PIN apb_paddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END apb_paddr[8]
  PIN apb_paddr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1465.440 1800.000 1466.040 ;
    END
  END apb_paddr[9]
  PIN apb_penable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1729.230 1796.000 1729.510 1800.000 ;
    END
  END apb_penable
  PIN apb_prdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END apb_prdata[0]
  PIN apb_prdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END apb_prdata[10]
  PIN apb_prdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 799.040 1800.000 799.640 ;
    END
  END apb_prdata[11]
  PIN apb_prdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 492.750 1796.000 493.030 1800.000 ;
    END
  END apb_prdata[12]
  PIN apb_prdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 945.240 1800.000 945.840 ;
    END
  END apb_prdata[13]
  PIN apb_prdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END apb_prdata[14]
  PIN apb_prdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 248.240 1800.000 248.840 ;
    END
  END apb_prdata[15]
  PIN apb_prdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 710.640 1800.000 711.240 ;
    END
  END apb_prdata[16]
  PIN apb_prdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1349.840 1800.000 1350.440 ;
    END
  END apb_prdata[17]
  PIN apb_prdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 1796.000 409.310 1800.000 ;
    END
  END apb_prdata[18]
  PIN apb_prdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END apb_prdata[19]
  PIN apb_prdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END apb_prdata[1]
  PIN apb_prdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END apb_prdata[20]
  PIN apb_prdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 1796.000 161.370 1800.000 ;
    END
  END apb_prdata[21]
  PIN apb_prdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1481.290 1796.000 1481.570 1800.000 ;
    END
  END apb_prdata[22]
  PIN apb_prdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 13.640 1800.000 14.240 ;
    END
  END apb_prdata[23]
  PIN apb_prdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END apb_prdata[24]
  PIN apb_prdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END apb_prdata[25]
  PIN apb_prdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END apb_prdata[26]
  PIN apb_prdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 930.670 1796.000 930.950 1800.000 ;
    END
  END apb_prdata[27]
  PIN apb_prdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END apb_prdata[28]
  PIN apb_prdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1593.990 0.000 1594.270 4.000 ;
    END
  END apb_prdata[29]
  PIN apb_prdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 884.040 1800.000 884.640 ;
    END
  END apb_prdata[2]
  PIN apb_prdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 1796.000 245.090 1800.000 ;
    END
  END apb_prdata[30]
  PIN apb_prdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END apb_prdata[31]
  PIN apb_prdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 795.430 1796.000 795.710 1800.000 ;
    END
  END apb_prdata[3]
  PIN apb_prdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END apb_prdata[4]
  PIN apb_prdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END apb_prdata[5]
  PIN apb_prdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 1796.000 1565.290 1800.000 ;
    END
  END apb_prdata[6]
  PIN apb_prdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END apb_prdata[7]
  PIN apb_prdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 1796.000 328.810 1800.000 ;
    END
  END apb_prdata[8]
  PIN apb_prdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END apb_prdata[9]
  PIN apb_pready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1700.040 1800.000 1700.640 ;
    END
  END apb_pready
  PIN apb_psel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END apb_psel
  PIN apb_pslverr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END apb_pslverr
  PIN apb_pwdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END apb_pwdata[0]
  PIN apb_pwdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 850.170 1796.000 850.450 1800.000 ;
    END
  END apb_pwdata[10]
  PIN apb_pwdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END apb_pwdata[11]
  PIN apb_pwdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1030.240 1800.000 1030.840 ;
    END
  END apb_pwdata[12]
  PIN apb_pwdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1619.750 1796.000 1620.030 1800.000 ;
    END
  END apb_pwdata[13]
  PIN apb_pwdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END apb_pwdata[14]
  PIN apb_pwdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 988.630 1796.000 988.910 1800.000 ;
    END
  END apb_pwdata[15]
  PIN apb_pwdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1796.000 1014.670 1800.000 ;
    END
  END apb_pwdata[16]
  PIN apb_pwdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1611.640 1800.000 1612.240 ;
    END
  END apb_pwdata[17]
  PIN apb_pwdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 740.690 1796.000 740.970 1800.000 ;
    END
  END apb_pwdata[18]
  PIN apb_pwdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END apb_pwdata[19]
  PIN apb_pwdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1203.640 1800.000 1204.240 ;
    END
  END apb_pwdata[1]
  PIN apb_pwdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END apb_pwdata[20]
  PIN apb_pwdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END apb_pwdata[21]
  PIN apb_pwdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END apb_pwdata[22]
  PIN apb_pwdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 1796.000 299.830 1800.000 ;
    END
  END apb_pwdata[23]
  PIN apb_pwdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 959.650 1796.000 959.930 1800.000 ;
    END
  END apb_pwdata[24]
  PIN apb_pwdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 972.440 1800.000 973.040 ;
    END
  END apb_pwdata[25]
  PIN apb_pwdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1455.530 1796.000 1455.810 1800.000 ;
    END
  END apb_pwdata[26]
  PIN apb_pwdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END apb_pwdata[27]
  PIN apb_pwdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 627.990 1796.000 628.270 1800.000 ;
    END
  END apb_pwdata[28]
  PIN apb_pwdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1796.000 1124.150 1800.000 ;
    END
  END apb_pwdata[29]
  PIN apb_pwdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 766.450 1796.000 766.730 1800.000 ;
    END
  END apb_pwdata[2]
  PIN apb_pwdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 1796.000 135.610 1800.000 ;
    END
  END apb_pwdata[30]
  PIN apb_pwdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END apb_pwdata[31]
  PIN apb_pwdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1060.840 1800.000 1061.440 ;
    END
  END apb_pwdata[3]
  PIN apb_pwdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1069.130 1796.000 1069.410 1800.000 ;
    END
  END apb_pwdata[4]
  PIN apb_pwdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1288.090 1796.000 1288.370 1800.000 ;
    END
  END apb_pwdata[5]
  PIN apb_pwdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END apb_pwdata[6]
  PIN apb_pwdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END apb_pwdata[7]
  PIN apb_pwdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END apb_pwdata[8]
  PIN apb_pwdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END apb_pwdata[9]
  PIN apb_pwrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END apb_pwrite
  PIN axi_aclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.721400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END axi_aclk
  PIN axi_araddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 391.040 1800.000 391.640 ;
    END
  END axi_araddr[0]
  PIN axi_araddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 479.440 1800.000 480.040 ;
    END
  END axi_araddr[10]
  PIN axi_araddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1727.240 1800.000 1727.840 ;
    END
  END axi_araddr[11]
  PIN axi_araddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 1796.000 1317.350 1800.000 ;
    END
  END axi_araddr[12]
  PIN axi_araddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 275.440 1800.000 276.040 ;
    END
  END axi_araddr[13]
  PIN axi_araddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 518.510 1796.000 518.790 1800.000 ;
    END
  END axi_araddr[14]
  PIN axi_araddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END axi_araddr[15]
  PIN axi_araddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END axi_araddr[16]
  PIN axi_araddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END axi_araddr[17]
  PIN axi_araddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END axi_araddr[18]
  PIN axi_araddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END axi_araddr[19]
  PIN axi_araddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END axi_araddr[1]
  PIN axi_araddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 652.840 1800.000 653.440 ;
    END
  END axi_araddr[20]
  PIN axi_araddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END axi_araddr[21]
  PIN axi_araddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END axi_araddr[22]
  PIN axi_araddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END axi_araddr[23]
  PIN axi_araddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END axi_araddr[24]
  PIN axi_araddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END axi_araddr[25]
  PIN axi_araddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 914.640 1800.000 915.240 ;
    END
  END axi_araddr[26]
  PIN axi_araddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1262.330 1796.000 1262.610 1800.000 ;
    END
  END axi_araddr[27]
  PIN axi_araddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 1796.000 190.350 1800.000 ;
    END
  END axi_araddr[28]
  PIN axi_araddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END axi_araddr[29]
  PIN axi_araddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END axi_araddr[2]
  PIN axi_araddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END axi_araddr[30]
  PIN axi_araddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END axi_araddr[31]
  PIN axi_araddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 821.190 1796.000 821.470 1800.000 ;
    END
  END axi_araddr[3]
  PIN axi_araddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END axi_araddr[4]
  PIN axi_araddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END axi_araddr[5]
  PIN axi_araddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1234.240 1800.000 1234.840 ;
    END
  END axi_araddr[6]
  PIN axi_araddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 159.840 1800.000 160.440 ;
    END
  END axi_araddr[7]
  PIN axi_araddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END axi_araddr[8]
  PIN axi_araddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1003.040 1800.000 1003.640 ;
    END
  END axi_araddr[9]
  PIN axi_aresetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END axi_aresetn
  PIN axi_arprot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1407.640 1800.000 1408.240 ;
    END
  END axi_arprot[0]
  PIN axi_arprot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END axi_arprot[1]
  PIN axi_arprot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 1796.000 1674.770 1800.000 ;
    END
  END axi_arprot[2]
  PIN axi_arready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END axi_arready
  PIN axi_arvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 187.040 1800.000 187.640 ;
    END
  END axi_arvalid
  PIN axi_awaddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END axi_awaddr[0]
  PIN axi_awaddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 448.840 1800.000 449.440 ;
    END
  END axi_awaddr[10]
  PIN axi_awaddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 1796.000 80.870 1800.000 ;
    END
  END axi_awaddr[11]
  PIN axi_awaddr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END axi_awaddr[12]
  PIN axi_awaddr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END axi_awaddr[13]
  PIN axi_awaddr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 547.490 1796.000 547.770 1800.000 ;
    END
  END axi_awaddr[14]
  PIN axi_awaddr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 625.640 1800.000 626.240 ;
    END
  END axi_awaddr[15]
  PIN axi_awaddr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1536.030 1796.000 1536.310 1800.000 ;
    END
  END axi_awaddr[16]
  PIN axi_awaddr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1648.730 1796.000 1649.010 1800.000 ;
    END
  END axi_awaddr[17]
  PIN axi_awaddr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END axi_awaddr[18]
  PIN axi_awaddr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1426.550 1796.000 1426.830 1800.000 ;
    END
  END axi_awaddr[19]
  PIN axi_awaddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 875.930 1796.000 876.210 1800.000 ;
    END
  END axi_awaddr[1]
  PIN axi_awaddr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END axi_awaddr[20]
  PIN axi_awaddr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1758.210 1796.000 1758.490 1800.000 ;
    END
  END axi_awaddr[21]
  PIN axi_awaddr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1796.000 1178.890 1800.000 ;
    END
  END axi_awaddr[22]
  PIN axi_awaddr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END axi_awaddr[23]
  PIN axi_awaddr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 656.970 1796.000 657.250 1800.000 ;
    END
  END axi_awaddr[24]
  PIN axi_awaddr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 683.440 1800.000 684.040 ;
    END
  END axi_awaddr[25]
  PIN axi_awaddr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 1796.000 51.890 1800.000 ;
    END
  END axi_awaddr[26]
  PIN axi_awaddr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END axi_awaddr[27]
  PIN axi_awaddr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 506.640 1800.000 507.240 ;
    END
  END axi_awaddr[28]
  PIN axi_awaddr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 71.440 1800.000 72.040 ;
    END
  END axi_awaddr[29]
  PIN axi_awaddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END axi_awaddr[2]
  PIN axi_awaddr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1669.440 1800.000 1670.040 ;
    END
  END axi_awaddr[30]
  PIN axi_awaddr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END axi_awaddr[31]
  PIN axi_awaddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END axi_awaddr[3]
  PIN axi_awaddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END axi_awaddr[4]
  PIN axi_awaddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END axi_awaddr[5]
  PIN axi_awaddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END axi_awaddr[6]
  PIN axi_awaddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END axi_awaddr[7]
  PIN axi_awaddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END axi_awaddr[8]
  PIN axi_awaddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END axi_awaddr[9]
  PIN axi_awprot[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END axi_awprot[0]
  PIN axi_awprot[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1176.440 1800.000 1177.040 ;
    END
  END axi_awprot[1]
  PIN axi_awprot[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END axi_awprot[2]
  PIN axi_awready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1581.040 1800.000 1581.640 ;
    END
  END axi_awready
  PIN axi_awvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END axi_awvalid
  PIN axi_bready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END axi_bready
  PIN axi_bresp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1642.240 1800.000 1642.840 ;
    END
  END axi_bresp[0]
  PIN axi_bresp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END axi_bresp[1]
  PIN axi_bvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END axi_bvalid
  PIN axi_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 1796.000 106.630 1800.000 ;
    END
  END axi_rdata[0]
  PIN axi_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END axi_rdata[10]
  PIN axi_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 129.240 1800.000 129.840 ;
    END
  END axi_rdata[11]
  PIN axi_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END axi_rdata[12]
  PIN axi_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1118.640 1800.000 1119.240 ;
    END
  END axi_rdata[13]
  PIN axi_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 354.290 1796.000 354.570 1800.000 ;
    END
  END axi_rdata[14]
  PIN axi_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 438.010 1796.000 438.290 1800.000 ;
    END
  END axi_rdata[15]
  PIN axi_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 383.270 1796.000 383.550 1800.000 ;
    END
  END axi_rdata[16]
  PIN axi_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END axi_rdata[17]
  PIN axi_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END axi_rdata[18]
  PIN axi_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 595.040 1800.000 595.640 ;
    END
  END axi_rdata[19]
  PIN axi_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END axi_rdata[1]
  PIN axi_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END axi_rdata[20]
  PIN axi_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1523.240 1800.000 1523.840 ;
    END
  END axi_rdata[21]
  PIN axi_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 685.950 1796.000 686.230 1800.000 ;
    END
  END axi_rdata[22]
  PIN axi_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END axi_rdata[23]
  PIN axi_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 768.440 1800.000 769.040 ;
    END
  END axi_rdata[24]
  PIN axi_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1496.040 1800.000 1496.640 ;
    END
  END axi_rdata[25]
  PIN axi_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END axi_rdata[26]
  PIN axi_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1088.040 1800.000 1088.640 ;
    END
  END axi_rdata[27]
  PIN axi_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 333.240 1800.000 333.840 ;
    END
  END axi_rdata[28]
  PIN axi_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END axi_rdata[29]
  PIN axi_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1757.840 1800.000 1758.440 ;
    END
  END axi_rdata[2]
  PIN axi_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 904.910 1796.000 905.190 1800.000 ;
    END
  END axi_rdata[30]
  PIN axi_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END axi_rdata[31]
  PIN axi_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END axi_rdata[3]
  PIN axi_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END axi_rdata[4]
  PIN axi_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 306.040 1800.000 306.640 ;
    END
  END axi_rdata[5]
  PIN axi_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END axi_rdata[6]
  PIN axi_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END axi_rdata[7]
  PIN axi_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END axi_rdata[8]
  PIN axi_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END axi_rdata[9]
  PIN axi_rready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 567.840 1800.000 568.440 ;
    END
  END axi_rready
  PIN axi_rresp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 1796.000 1703.750 1800.000 ;
    END
  END axi_rresp[0]
  PIN axi_rresp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1380.440 1800.000 1381.040 ;
    END
  END axi_rresp[1]
  PIN axi_rvalid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END axi_rvalid
  PIN axi_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END axi_wdata[0]
  PIN axi_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 826.240 1800.000 826.840 ;
    END
  END axi_wdata[10]
  PIN axi_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END axi_wdata[11]
  PIN axi_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1438.240 1800.000 1438.840 ;
    END
  END axi_wdata[12]
  PIN axi_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1590.770 1796.000 1591.050 1800.000 ;
    END
  END axi_wdata[13]
  PIN axi_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 44.240 1800.000 44.840 ;
    END
  END axi_wdata[14]
  PIN axi_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 1796.000 1510.550 1800.000 ;
    END
  END axi_wdata[15]
  PIN axi_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END axi_wdata[16]
  PIN axi_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END axi_wdata[17]
  PIN axi_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END axi_wdata[18]
  PIN axi_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END axi_wdata[19]
  PIN axi_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END axi_wdata[1]
  PIN axi_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END axi_wdata[20]
  PIN axi_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 1796.000 26.130 1800.000 ;
    END
  END axi_wdata[21]
  PIN axi_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END axi_wdata[22]
  PIN axi_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END axi_wdata[23]
  PIN axi_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END axi_wdata[24]
  PIN axi_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END axi_wdata[25]
  PIN axi_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1796.000 1098.390 1800.000 ;
    END
  END axi_wdata[26]
  PIN axi_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 711.710 1796.000 711.990 1800.000 ;
    END
  END axi_wdata[27]
  PIN axi_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END axi_wdata[28]
  PIN axi_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1371.810 1796.000 1372.090 1800.000 ;
    END
  END axi_wdata[29]
  PIN axi_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 421.640 1800.000 422.240 ;
    END
  END axi_wdata[2]
  PIN axi_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END axi_wdata[30]
  PIN axi_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1322.640 1800.000 1323.240 ;
    END
  END axi_wdata[31]
  PIN axi_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END axi_wdata[3]
  PIN axi_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END axi_wdata[4]
  PIN axi_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END axi_wdata[5]
  PIN axi_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1261.440 1800.000 1262.040 ;
    END
  END axi_wdata[6]
  PIN axi_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END axi_wdata[7]
  PIN axi_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1796.000 1233.630 1800.000 ;
    END
  END axi_wdata[8]
  PIN axi_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1207.590 1796.000 1207.870 1800.000 ;
    END
  END axi_wdata[9]
  PIN axi_wready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1771.440 4.000 1772.040 ;
    END
  END axi_wready
  PIN axi_wstrb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1796.000 270.850 1800.000 ;
    END
  END axi_wstrb[0]
  PIN axi_wstrb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END axi_wstrb[1]
  PIN axi_wstrb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END axi_wstrb[2]
  PIN axi_wstrb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END axi_wstrb[3]
  PIN axi_wvalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 1796.000 856.840 1800.000 857.440 ;
    END
  END axi_wvalid
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1794.460 1787.125 ;
      LAYER met1 ;
        RECT 0.070 8.200 1795.310 1787.280 ;
      LAYER met2 ;
        RECT 0.100 1795.720 25.570 1799.125 ;
        RECT 26.410 1795.720 51.330 1799.125 ;
        RECT 52.170 1795.720 80.310 1799.125 ;
        RECT 81.150 1795.720 106.070 1799.125 ;
        RECT 106.910 1795.720 135.050 1799.125 ;
        RECT 135.890 1795.720 160.810 1799.125 ;
        RECT 161.650 1795.720 189.790 1799.125 ;
        RECT 190.630 1795.720 215.550 1799.125 ;
        RECT 216.390 1795.720 244.530 1799.125 ;
        RECT 245.370 1795.720 270.290 1799.125 ;
        RECT 271.130 1795.720 299.270 1799.125 ;
        RECT 300.110 1795.720 328.250 1799.125 ;
        RECT 329.090 1795.720 354.010 1799.125 ;
        RECT 354.850 1795.720 382.990 1799.125 ;
        RECT 383.830 1795.720 408.750 1799.125 ;
        RECT 409.590 1795.720 437.730 1799.125 ;
        RECT 438.570 1795.720 463.490 1799.125 ;
        RECT 464.330 1795.720 492.470 1799.125 ;
        RECT 493.310 1795.720 518.230 1799.125 ;
        RECT 519.070 1795.720 547.210 1799.125 ;
        RECT 548.050 1795.720 572.970 1799.125 ;
        RECT 573.810 1795.720 601.950 1799.125 ;
        RECT 602.790 1795.720 627.710 1799.125 ;
        RECT 628.550 1795.720 656.690 1799.125 ;
        RECT 657.530 1795.720 685.670 1799.125 ;
        RECT 686.510 1795.720 711.430 1799.125 ;
        RECT 712.270 1795.720 740.410 1799.125 ;
        RECT 741.250 1795.720 766.170 1799.125 ;
        RECT 767.010 1795.720 795.150 1799.125 ;
        RECT 795.990 1795.720 820.910 1799.125 ;
        RECT 821.750 1795.720 849.890 1799.125 ;
        RECT 850.730 1795.720 875.650 1799.125 ;
        RECT 876.490 1795.720 904.630 1799.125 ;
        RECT 905.470 1795.720 930.390 1799.125 ;
        RECT 931.230 1795.720 959.370 1799.125 ;
        RECT 960.210 1795.720 988.350 1799.125 ;
        RECT 989.190 1795.720 1014.110 1799.125 ;
        RECT 1014.950 1795.720 1043.090 1799.125 ;
        RECT 1043.930 1795.720 1068.850 1799.125 ;
        RECT 1069.690 1795.720 1097.830 1799.125 ;
        RECT 1098.670 1795.720 1123.590 1799.125 ;
        RECT 1124.430 1795.720 1152.570 1799.125 ;
        RECT 1153.410 1795.720 1178.330 1799.125 ;
        RECT 1179.170 1795.720 1207.310 1799.125 ;
        RECT 1208.150 1795.720 1233.070 1799.125 ;
        RECT 1233.910 1795.720 1262.050 1799.125 ;
        RECT 1262.890 1795.720 1287.810 1799.125 ;
        RECT 1288.650 1795.720 1316.790 1799.125 ;
        RECT 1317.630 1795.720 1345.770 1799.125 ;
        RECT 1346.610 1795.720 1371.530 1799.125 ;
        RECT 1372.370 1795.720 1400.510 1799.125 ;
        RECT 1401.350 1795.720 1426.270 1799.125 ;
        RECT 1427.110 1795.720 1455.250 1799.125 ;
        RECT 1456.090 1795.720 1481.010 1799.125 ;
        RECT 1481.850 1795.720 1509.990 1799.125 ;
        RECT 1510.830 1795.720 1535.750 1799.125 ;
        RECT 1536.590 1795.720 1564.730 1799.125 ;
        RECT 1565.570 1795.720 1590.490 1799.125 ;
        RECT 1591.330 1795.720 1619.470 1799.125 ;
        RECT 1620.310 1795.720 1648.450 1799.125 ;
        RECT 1649.290 1795.720 1674.210 1799.125 ;
        RECT 1675.050 1795.720 1703.190 1799.125 ;
        RECT 1704.030 1795.720 1728.950 1799.125 ;
        RECT 1729.790 1795.720 1757.930 1799.125 ;
        RECT 1758.770 1795.720 1783.690 1799.125 ;
        RECT 1784.530 1795.720 1795.290 1799.125 ;
        RECT 0.100 4.280 1795.290 1795.720 ;
        RECT 0.650 3.670 25.570 4.280 ;
        RECT 26.410 3.670 54.550 4.280 ;
        RECT 55.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 109.290 4.280 ;
        RECT 110.130 3.670 135.050 4.280 ;
        RECT 135.890 3.670 164.030 4.280 ;
        RECT 164.870 3.670 189.790 4.280 ;
        RECT 190.630 3.670 218.770 4.280 ;
        RECT 219.610 3.670 244.530 4.280 ;
        RECT 245.370 3.670 273.510 4.280 ;
        RECT 274.350 3.670 299.270 4.280 ;
        RECT 300.110 3.670 328.250 4.280 ;
        RECT 329.090 3.670 357.230 4.280 ;
        RECT 358.070 3.670 382.990 4.280 ;
        RECT 383.830 3.670 411.970 4.280 ;
        RECT 412.810 3.670 437.730 4.280 ;
        RECT 438.570 3.670 466.710 4.280 ;
        RECT 467.550 3.670 492.470 4.280 ;
        RECT 493.310 3.670 521.450 4.280 ;
        RECT 522.290 3.670 547.210 4.280 ;
        RECT 548.050 3.670 576.190 4.280 ;
        RECT 577.030 3.670 601.950 4.280 ;
        RECT 602.790 3.670 630.930 4.280 ;
        RECT 631.770 3.670 656.690 4.280 ;
        RECT 657.530 3.670 685.670 4.280 ;
        RECT 686.510 3.670 714.650 4.280 ;
        RECT 715.490 3.670 740.410 4.280 ;
        RECT 741.250 3.670 769.390 4.280 ;
        RECT 770.230 3.670 795.150 4.280 ;
        RECT 795.990 3.670 824.130 4.280 ;
        RECT 824.970 3.670 849.890 4.280 ;
        RECT 850.730 3.670 878.870 4.280 ;
        RECT 879.710 3.670 904.630 4.280 ;
        RECT 905.470 3.670 933.610 4.280 ;
        RECT 934.450 3.670 959.370 4.280 ;
        RECT 960.210 3.670 988.350 4.280 ;
        RECT 989.190 3.670 1017.330 4.280 ;
        RECT 1018.170 3.670 1043.090 4.280 ;
        RECT 1043.930 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1126.810 4.280 ;
        RECT 1127.650 3.670 1152.570 4.280 ;
        RECT 1153.410 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1207.310 4.280 ;
        RECT 1208.150 3.670 1236.290 4.280 ;
        RECT 1237.130 3.670 1262.050 4.280 ;
        RECT 1262.890 3.670 1291.030 4.280 ;
        RECT 1291.870 3.670 1316.790 4.280 ;
        RECT 1317.630 3.670 1345.770 4.280 ;
        RECT 1346.610 3.670 1374.750 4.280 ;
        RECT 1375.590 3.670 1400.510 4.280 ;
        RECT 1401.350 3.670 1429.490 4.280 ;
        RECT 1430.330 3.670 1455.250 4.280 ;
        RECT 1456.090 3.670 1484.230 4.280 ;
        RECT 1485.070 3.670 1509.990 4.280 ;
        RECT 1510.830 3.670 1538.970 4.280 ;
        RECT 1539.810 3.670 1564.730 4.280 ;
        RECT 1565.570 3.670 1593.710 4.280 ;
        RECT 1594.550 3.670 1619.470 4.280 ;
        RECT 1620.310 3.670 1648.450 4.280 ;
        RECT 1649.290 3.670 1677.430 4.280 ;
        RECT 1678.270 3.670 1703.190 4.280 ;
        RECT 1704.030 3.670 1732.170 4.280 ;
        RECT 1733.010 3.670 1757.930 4.280 ;
        RECT 1758.770 3.670 1786.910 4.280 ;
        RECT 1787.750 3.670 1795.290 4.280 ;
      LAYER met3 ;
        RECT 4.400 1798.240 1796.000 1799.105 ;
        RECT 3.990 1786.040 1796.000 1798.240 ;
        RECT 3.990 1784.640 1795.600 1786.040 ;
        RECT 3.990 1772.440 1796.000 1784.640 ;
        RECT 4.400 1771.040 1796.000 1772.440 ;
        RECT 3.990 1758.840 1796.000 1771.040 ;
        RECT 3.990 1757.440 1795.600 1758.840 ;
        RECT 3.990 1741.840 1796.000 1757.440 ;
        RECT 4.400 1740.440 1796.000 1741.840 ;
        RECT 3.990 1728.240 1796.000 1740.440 ;
        RECT 3.990 1726.840 1795.600 1728.240 ;
        RECT 3.990 1711.240 1796.000 1726.840 ;
        RECT 4.400 1709.840 1796.000 1711.240 ;
        RECT 3.990 1701.040 1796.000 1709.840 ;
        RECT 3.990 1699.640 1795.600 1701.040 ;
        RECT 3.990 1684.040 1796.000 1699.640 ;
        RECT 4.400 1682.640 1796.000 1684.040 ;
        RECT 3.990 1670.440 1796.000 1682.640 ;
        RECT 3.990 1669.040 1795.600 1670.440 ;
        RECT 3.990 1653.440 1796.000 1669.040 ;
        RECT 4.400 1652.040 1796.000 1653.440 ;
        RECT 3.990 1643.240 1796.000 1652.040 ;
        RECT 3.990 1641.840 1795.600 1643.240 ;
        RECT 3.990 1626.240 1796.000 1641.840 ;
        RECT 4.400 1624.840 1796.000 1626.240 ;
        RECT 3.990 1612.640 1796.000 1624.840 ;
        RECT 3.990 1611.240 1795.600 1612.640 ;
        RECT 3.990 1595.640 1796.000 1611.240 ;
        RECT 4.400 1594.240 1796.000 1595.640 ;
        RECT 3.990 1582.040 1796.000 1594.240 ;
        RECT 3.990 1580.640 1795.600 1582.040 ;
        RECT 3.990 1568.440 1796.000 1580.640 ;
        RECT 4.400 1567.040 1796.000 1568.440 ;
        RECT 3.990 1554.840 1796.000 1567.040 ;
        RECT 3.990 1553.440 1795.600 1554.840 ;
        RECT 3.990 1537.840 1796.000 1553.440 ;
        RECT 4.400 1536.440 1796.000 1537.840 ;
        RECT 3.990 1524.240 1796.000 1536.440 ;
        RECT 3.990 1522.840 1795.600 1524.240 ;
        RECT 3.990 1510.640 1796.000 1522.840 ;
        RECT 4.400 1509.240 1796.000 1510.640 ;
        RECT 3.990 1497.040 1796.000 1509.240 ;
        RECT 3.990 1495.640 1795.600 1497.040 ;
        RECT 3.990 1480.040 1796.000 1495.640 ;
        RECT 4.400 1478.640 1796.000 1480.040 ;
        RECT 3.990 1466.440 1796.000 1478.640 ;
        RECT 3.990 1465.040 1795.600 1466.440 ;
        RECT 3.990 1452.840 1796.000 1465.040 ;
        RECT 4.400 1451.440 1796.000 1452.840 ;
        RECT 3.990 1439.240 1796.000 1451.440 ;
        RECT 3.990 1437.840 1795.600 1439.240 ;
        RECT 3.990 1422.240 1796.000 1437.840 ;
        RECT 4.400 1420.840 1796.000 1422.240 ;
        RECT 3.990 1408.640 1796.000 1420.840 ;
        RECT 3.990 1407.240 1795.600 1408.640 ;
        RECT 3.990 1391.640 1796.000 1407.240 ;
        RECT 4.400 1390.240 1796.000 1391.640 ;
        RECT 3.990 1381.440 1796.000 1390.240 ;
        RECT 3.990 1380.040 1795.600 1381.440 ;
        RECT 3.990 1364.440 1796.000 1380.040 ;
        RECT 4.400 1363.040 1796.000 1364.440 ;
        RECT 3.990 1350.840 1796.000 1363.040 ;
        RECT 3.990 1349.440 1795.600 1350.840 ;
        RECT 3.990 1333.840 1796.000 1349.440 ;
        RECT 4.400 1332.440 1796.000 1333.840 ;
        RECT 3.990 1323.640 1796.000 1332.440 ;
        RECT 3.990 1322.240 1795.600 1323.640 ;
        RECT 3.990 1306.640 1796.000 1322.240 ;
        RECT 4.400 1305.240 1796.000 1306.640 ;
        RECT 3.990 1293.040 1796.000 1305.240 ;
        RECT 3.990 1291.640 1795.600 1293.040 ;
        RECT 3.990 1276.040 1796.000 1291.640 ;
        RECT 4.400 1274.640 1796.000 1276.040 ;
        RECT 3.990 1262.440 1796.000 1274.640 ;
        RECT 3.990 1261.040 1795.600 1262.440 ;
        RECT 3.990 1248.840 1796.000 1261.040 ;
        RECT 4.400 1247.440 1796.000 1248.840 ;
        RECT 3.990 1235.240 1796.000 1247.440 ;
        RECT 3.990 1233.840 1795.600 1235.240 ;
        RECT 3.990 1218.240 1796.000 1233.840 ;
        RECT 4.400 1216.840 1796.000 1218.240 ;
        RECT 3.990 1204.640 1796.000 1216.840 ;
        RECT 3.990 1203.240 1795.600 1204.640 ;
        RECT 3.990 1191.040 1796.000 1203.240 ;
        RECT 4.400 1189.640 1796.000 1191.040 ;
        RECT 3.990 1177.440 1796.000 1189.640 ;
        RECT 3.990 1176.040 1795.600 1177.440 ;
        RECT 3.990 1160.440 1796.000 1176.040 ;
        RECT 4.400 1159.040 1796.000 1160.440 ;
        RECT 3.990 1146.840 1796.000 1159.040 ;
        RECT 3.990 1145.440 1795.600 1146.840 ;
        RECT 3.990 1133.240 1796.000 1145.440 ;
        RECT 4.400 1131.840 1796.000 1133.240 ;
        RECT 3.990 1119.640 1796.000 1131.840 ;
        RECT 3.990 1118.240 1795.600 1119.640 ;
        RECT 3.990 1102.640 1796.000 1118.240 ;
        RECT 4.400 1101.240 1796.000 1102.640 ;
        RECT 3.990 1089.040 1796.000 1101.240 ;
        RECT 3.990 1087.640 1795.600 1089.040 ;
        RECT 3.990 1075.440 1796.000 1087.640 ;
        RECT 4.400 1074.040 1796.000 1075.440 ;
        RECT 3.990 1061.840 1796.000 1074.040 ;
        RECT 3.990 1060.440 1795.600 1061.840 ;
        RECT 3.990 1044.840 1796.000 1060.440 ;
        RECT 4.400 1043.440 1796.000 1044.840 ;
        RECT 3.990 1031.240 1796.000 1043.440 ;
        RECT 3.990 1029.840 1795.600 1031.240 ;
        RECT 3.990 1014.240 1796.000 1029.840 ;
        RECT 4.400 1012.840 1796.000 1014.240 ;
        RECT 3.990 1004.040 1796.000 1012.840 ;
        RECT 3.990 1002.640 1795.600 1004.040 ;
        RECT 3.990 987.040 1796.000 1002.640 ;
        RECT 4.400 985.640 1796.000 987.040 ;
        RECT 3.990 973.440 1796.000 985.640 ;
        RECT 3.990 972.040 1795.600 973.440 ;
        RECT 3.990 956.440 1796.000 972.040 ;
        RECT 4.400 955.040 1796.000 956.440 ;
        RECT 3.990 946.240 1796.000 955.040 ;
        RECT 3.990 944.840 1795.600 946.240 ;
        RECT 3.990 929.240 1796.000 944.840 ;
        RECT 4.400 927.840 1796.000 929.240 ;
        RECT 3.990 915.640 1796.000 927.840 ;
        RECT 3.990 914.240 1795.600 915.640 ;
        RECT 3.990 898.640 1796.000 914.240 ;
        RECT 4.400 897.240 1796.000 898.640 ;
        RECT 3.990 885.040 1796.000 897.240 ;
        RECT 3.990 883.640 1795.600 885.040 ;
        RECT 3.990 871.440 1796.000 883.640 ;
        RECT 4.400 870.040 1796.000 871.440 ;
        RECT 3.990 857.840 1796.000 870.040 ;
        RECT 3.990 856.440 1795.600 857.840 ;
        RECT 3.990 840.840 1796.000 856.440 ;
        RECT 4.400 839.440 1796.000 840.840 ;
        RECT 3.990 827.240 1796.000 839.440 ;
        RECT 3.990 825.840 1795.600 827.240 ;
        RECT 3.990 813.640 1796.000 825.840 ;
        RECT 4.400 812.240 1796.000 813.640 ;
        RECT 3.990 800.040 1796.000 812.240 ;
        RECT 3.990 798.640 1795.600 800.040 ;
        RECT 3.990 783.040 1796.000 798.640 ;
        RECT 4.400 781.640 1796.000 783.040 ;
        RECT 3.990 769.440 1796.000 781.640 ;
        RECT 3.990 768.040 1795.600 769.440 ;
        RECT 3.990 755.840 1796.000 768.040 ;
        RECT 4.400 754.440 1796.000 755.840 ;
        RECT 3.990 742.240 1796.000 754.440 ;
        RECT 3.990 740.840 1795.600 742.240 ;
        RECT 3.990 725.240 1796.000 740.840 ;
        RECT 4.400 723.840 1796.000 725.240 ;
        RECT 3.990 711.640 1796.000 723.840 ;
        RECT 3.990 710.240 1795.600 711.640 ;
        RECT 3.990 694.640 1796.000 710.240 ;
        RECT 4.400 693.240 1796.000 694.640 ;
        RECT 3.990 684.440 1796.000 693.240 ;
        RECT 3.990 683.040 1795.600 684.440 ;
        RECT 3.990 667.440 1796.000 683.040 ;
        RECT 4.400 666.040 1796.000 667.440 ;
        RECT 3.990 653.840 1796.000 666.040 ;
        RECT 3.990 652.440 1795.600 653.840 ;
        RECT 3.990 636.840 1796.000 652.440 ;
        RECT 4.400 635.440 1796.000 636.840 ;
        RECT 3.990 626.640 1796.000 635.440 ;
        RECT 3.990 625.240 1795.600 626.640 ;
        RECT 3.990 609.640 1796.000 625.240 ;
        RECT 4.400 608.240 1796.000 609.640 ;
        RECT 3.990 596.040 1796.000 608.240 ;
        RECT 3.990 594.640 1795.600 596.040 ;
        RECT 3.990 579.040 1796.000 594.640 ;
        RECT 4.400 577.640 1796.000 579.040 ;
        RECT 3.990 568.840 1796.000 577.640 ;
        RECT 3.990 567.440 1795.600 568.840 ;
        RECT 3.990 551.840 1796.000 567.440 ;
        RECT 4.400 550.440 1796.000 551.840 ;
        RECT 3.990 538.240 1796.000 550.440 ;
        RECT 3.990 536.840 1795.600 538.240 ;
        RECT 3.990 521.240 1796.000 536.840 ;
        RECT 4.400 519.840 1796.000 521.240 ;
        RECT 3.990 507.640 1796.000 519.840 ;
        RECT 3.990 506.240 1795.600 507.640 ;
        RECT 3.990 494.040 1796.000 506.240 ;
        RECT 4.400 492.640 1796.000 494.040 ;
        RECT 3.990 480.440 1796.000 492.640 ;
        RECT 3.990 479.040 1795.600 480.440 ;
        RECT 3.990 463.440 1796.000 479.040 ;
        RECT 4.400 462.040 1796.000 463.440 ;
        RECT 3.990 449.840 1796.000 462.040 ;
        RECT 3.990 448.440 1795.600 449.840 ;
        RECT 3.990 436.240 1796.000 448.440 ;
        RECT 4.400 434.840 1796.000 436.240 ;
        RECT 3.990 422.640 1796.000 434.840 ;
        RECT 3.990 421.240 1795.600 422.640 ;
        RECT 3.990 405.640 1796.000 421.240 ;
        RECT 4.400 404.240 1796.000 405.640 ;
        RECT 3.990 392.040 1796.000 404.240 ;
        RECT 3.990 390.640 1795.600 392.040 ;
        RECT 3.990 378.440 1796.000 390.640 ;
        RECT 4.400 377.040 1796.000 378.440 ;
        RECT 3.990 364.840 1796.000 377.040 ;
        RECT 3.990 363.440 1795.600 364.840 ;
        RECT 3.990 347.840 1796.000 363.440 ;
        RECT 4.400 346.440 1796.000 347.840 ;
        RECT 3.990 334.240 1796.000 346.440 ;
        RECT 3.990 332.840 1795.600 334.240 ;
        RECT 3.990 317.240 1796.000 332.840 ;
        RECT 4.400 315.840 1796.000 317.240 ;
        RECT 3.990 307.040 1796.000 315.840 ;
        RECT 3.990 305.640 1795.600 307.040 ;
        RECT 3.990 290.040 1796.000 305.640 ;
        RECT 4.400 288.640 1796.000 290.040 ;
        RECT 3.990 276.440 1796.000 288.640 ;
        RECT 3.990 275.040 1795.600 276.440 ;
        RECT 3.990 259.440 1796.000 275.040 ;
        RECT 4.400 258.040 1796.000 259.440 ;
        RECT 3.990 249.240 1796.000 258.040 ;
        RECT 3.990 247.840 1795.600 249.240 ;
        RECT 3.990 232.240 1796.000 247.840 ;
        RECT 4.400 230.840 1796.000 232.240 ;
        RECT 3.990 218.640 1796.000 230.840 ;
        RECT 3.990 217.240 1795.600 218.640 ;
        RECT 3.990 201.640 1796.000 217.240 ;
        RECT 4.400 200.240 1796.000 201.640 ;
        RECT 3.990 188.040 1796.000 200.240 ;
        RECT 3.990 186.640 1795.600 188.040 ;
        RECT 3.990 174.440 1796.000 186.640 ;
        RECT 4.400 173.040 1796.000 174.440 ;
        RECT 3.990 160.840 1796.000 173.040 ;
        RECT 3.990 159.440 1795.600 160.840 ;
        RECT 3.990 143.840 1796.000 159.440 ;
        RECT 4.400 142.440 1796.000 143.840 ;
        RECT 3.990 130.240 1796.000 142.440 ;
        RECT 3.990 128.840 1795.600 130.240 ;
        RECT 3.990 116.640 1796.000 128.840 ;
        RECT 4.400 115.240 1796.000 116.640 ;
        RECT 3.990 103.040 1796.000 115.240 ;
        RECT 3.990 101.640 1795.600 103.040 ;
        RECT 3.990 86.040 1796.000 101.640 ;
        RECT 4.400 84.640 1796.000 86.040 ;
        RECT 3.990 72.440 1796.000 84.640 ;
        RECT 3.990 71.040 1795.600 72.440 ;
        RECT 3.990 58.840 1796.000 71.040 ;
        RECT 4.400 57.440 1796.000 58.840 ;
        RECT 3.990 45.240 1796.000 57.440 ;
        RECT 3.990 43.840 1795.600 45.240 ;
        RECT 3.990 28.240 1796.000 43.840 ;
        RECT 4.400 26.840 1796.000 28.240 ;
        RECT 3.990 14.640 1796.000 26.840 ;
        RECT 3.990 13.240 1795.600 14.640 ;
        RECT 3.990 10.715 1796.000 13.240 ;
      LAYER met4 ;
        RECT 17.775 172.215 164.920 1622.305 ;
        RECT 167.320 172.215 168.220 1622.305 ;
        RECT 170.620 172.215 318.520 1622.305 ;
        RECT 320.920 172.215 321.820 1622.305 ;
        RECT 324.220 172.215 472.120 1622.305 ;
        RECT 474.520 172.215 475.420 1622.305 ;
        RECT 477.820 172.215 625.720 1622.305 ;
        RECT 628.120 172.215 629.020 1622.305 ;
        RECT 631.420 172.215 779.320 1622.305 ;
        RECT 781.720 172.215 782.620 1622.305 ;
        RECT 785.020 172.215 932.920 1622.305 ;
        RECT 935.320 172.215 936.220 1622.305 ;
        RECT 938.620 172.215 1086.520 1622.305 ;
        RECT 1088.920 172.215 1089.820 1622.305 ;
        RECT 1092.220 172.215 1240.120 1622.305 ;
        RECT 1242.520 172.215 1243.420 1622.305 ;
        RECT 1245.820 172.215 1393.720 1622.305 ;
        RECT 1396.120 172.215 1397.020 1622.305 ;
        RECT 1399.420 172.215 1448.705 1622.305 ;
  END
END axi_apb_bridge
END LIBRARY

